
module Chenillard_sys (
	clk_clk,
	reset_reset_n,
	leds_external_connection_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[7:0]	leds_external_connection_export;
endmodule
