
module Chenillard_sys (
	button_external_connection_export,
	clk_clk,
	leds_external_connection_export,
	reset_reset_n);	

	input		button_external_connection_export;
	input		clk_clk;
	output	[7:0]	leds_external_connection_export;
	input		reset_reset_n;
endmodule
